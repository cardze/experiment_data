library verilog;
use verilog.vl_types.all;
entity tes_013_vlg_vec_tst is
end tes_013_vlg_vec_tst;
