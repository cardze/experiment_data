library verilog;
use verilog.vl_types.all;
entity test_not_A_and_b_vlg_check_tst is
    port(
        result          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end test_not_A_and_b_vlg_check_tst;
