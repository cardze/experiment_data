library verilog;
use verilog.vl_types.all;
entity tes_013 is
    port(
        input_A         : in     vl_logic;
        input_B         : in     vl_logic;
        result          : out    vl_logic
    );
end tes_013;
