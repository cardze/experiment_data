library verilog;
use verilog.vl_types.all;
entity test_not_A_and_b_vlg_vec_tst is
end test_not_A_and_b_vlg_vec_tst;
