library verilog;
use verilog.vl_types.all;
entity test_ab_and_bc_vlg_vec_tst is
end test_ab_and_bc_vlg_vec_tst;
